library ieee;
use ieee.std_logic_1164.all;

ENTITY Decode IS
PORT(A,B,C,D,E: IN BIT;
S0,S1,S2,S3,S4,S5,S6 : OUT BIT);
END;
ARCHITECTURE behav OF Decode IS
BEGIN
S0 <= NOT(E) OR (NOT(A) AND NOT(B) AND NOT(C) AND D) OR (NOT(A) AND B AND NOT(C) AND NOT(D)) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S1 <= NOT(E) OR (NOT(A) AND B AND NOT(C) AND D) OR (NOT(A) AND B AND C AND NOT(D)) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S2 <= NOT(E) OR (NOT(A) AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S3 <= NOT(E) OR (NOT(A) AND NOT(B) AND NOT(C) AND D) OR (NOT(A) AND B AND NOT(C) AND NOT(D)) OR (NOT(A) AND B AND C AND D) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S4 <= NOT(E) OR (NOT(A) AND D) OR (NOT(A) AND B AND NOT(C)) OR (NOT(B) AND NOT(C) AND D) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S5 <= NOT(E) OR (NOT(A) AND NOT(B) AND C) OR (NOT(A) AND NOT(B) AND D) OR (NOT(A) AND C AND D) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
S6 <= NOT(E) OR (NOT(A) AND NOT(B) AND NOT(C)) OR (NOT(A) AND B AND C AND D) OR (A AND NOT(B) AND C AND NOT(D)) OR (A AND NOT(B) AND C AND D) OR (A AND B AND NOT(C) AND NOT(D)) OR (A AND B AND NOT(C) AND D) OR (A AND B AND C AND NOT(D)) OR (A AND B AND C AND D);
END;
